module shift_add_multiplier (
    input logic clk, rst,
    input logic[7:0] a,
    input logic[7:0] b,

    output logic[15:0] result,
    output logic d_end
);

    shift_register A (

    );

    shift_register B (

    );

    shift_register Q (

    );

    counter count (

    );

endmodule