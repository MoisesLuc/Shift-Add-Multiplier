module shift_add_multiplier (
    input logic clk, rst,
    input logic[7:0] a,
    input logic[7:0] b,

    output logic[15:0] result,
    output logic d_end
);

endmodule